
module lls #(
    parameter OPERAND_WIDTH = 4
) (
    input logic [OPERAND_WIDTH-1:0] x,
    input logic [$clog2(OPERAND_WIDTH)-1:0] y,
    output logic [OPERAND_WIDTH-1:0] z
);


assign z = x<<y;
    
endmodule;

// module lls #(
//     parameter OPERAND_WIDTH = 4
// ) (
//     input  logic [      OPERAND_WIDTH-1 : 0] x,
//     input  logic [$clog2(OPERAND_WIDTH)-1:0] y,
//     output logic [        OPERAND_WIDTH-1:0] z
// );

//   assign z = x << y;

// endmodule
// ;

// module and_gate(
//     input logic x,
//     input logic y,
//     output logic z
// );

//     assign z = x & y;
// endmodule;

module and_gate (
    input  logic x,
    input  logic y,
    output logic z
);
// 
  assign z = x & y;
// 
endmodule;

